`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/17/2017 05:35:13 PM
// Design Name: 
// Module Name: CIRCUIT1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module CIRCUIT5(a, b, c, x, z);
    
    input [63:0] a, b, c;
    output [31:0] x, z;
    
    reg [63:0] greg, hreg;
    
    wire [63:0] d, e, f, g, h; 
    wire dLTe, dEQe;
    wire [63:0] xrin, zrin;
    
endmodule