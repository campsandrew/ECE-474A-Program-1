`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Names: Andrew Camps, Jason Tran
// Create Date: 09/17/2017 05:35:13 PM
// Module Name: CIRCUIT1
//////////////////////////////////////////////////////////////////////////////////


module CIRCUIT4(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, final);
    
    input [7:0] a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p;
    output [31:0] final;
    
    wire [31:0] t1, t2, t3, t4, t5, t6, t7, t8, t9, t10, t11, t12, t13, t14;
    
    


endmodule